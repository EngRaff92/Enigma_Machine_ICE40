//! Configuration selector for Enigma 
//!

module config_selector(
    // Input Ports
    // Output Ports
);
endmodule // config_selector