module apb_master #(
    //! parameters
) (
    //! port_list
);
    
endmodule // apb_master