module enigma #(
    //
) (
    //
);
    
endmodule // enigma